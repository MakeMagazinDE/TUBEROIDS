-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ASTEROIDS_VEC_ROM_2 is
  port (
    CLK         : in    std_logic;
    ADDR        : in    std_logic_vector(10 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ASTEROIDS_VEC_ROM_2 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INITP_00 : string;
  attribute INITP_01 : string;
  attribute INITP_02 : string;
  attribute INITP_03 : string;
  attribute INITP_04 : string;
  attribute INITP_05 : string;
  attribute INITP_06 : string;
  attribute INITP_07 : string;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S9
    --pragma translate_off
    generic (
      INITP_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INITP_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";

      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (7 downto 0);
      DOP   : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (10 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (7 downto 0);
      DIP   : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(10 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(10 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "FE0AFF08FE0EF80FFA0E038051804FCE4F9E4F6A4F3A4F064ED24E9E4E847680";
    attribute INIT_01 of inst : label is "C89FC896C88DC884C87BC872C869C860C857C84EC84507805580FB08FA0AF80B";
    attribute INIT_02 of inst : label is "C92FC926C91DC914C90BC902C8F9C8F0C8E7C8DEC8D5C8CCC8C3C8BAC8B1C8A8";
    attribute INIT_03 of inst : label is "C99DC997C993C98DC987C981C97BC975C96FC969C965C95CC953C94AC941C938";
    attribute INIT_04 of inst : label is "76A04300D00072004380770055C0730055C076004380C9BBC9B5C9AFC9A9C9A3";
    attribute INIT_05 of inst : label is "D00070405200762056C07370548077204280D000714043E07690565073405520";
    attribute INIT_06 of inst : label is "43E074F05760736050F077E04100D00074205200759057207380504077A041C0";
    attribute INIT_07 of inst : label is "577072C0522076005440D00075C043A0744057807320519076005020D0007500";
    attribute INIT_08 of inst : label is "530077804600D000770042A0712057407250529077E04540D000768043207080";
    attribute INIT_09 of inst : label is "4720D00077E041407250569071205340770046A0D0007780420071C0570071C0";
    attribute INIT_0A of inst : label is "76005420732055907440538075C047A0D0007600504072C05620708053707680";
    attribute INIT_0B of inst : label is "738054407590532074205600D00077E04500736054F074F05360750047E0D000";
    attribute INIT_0C of inst : label is "76905250714047E0D0007720468073705080762052C070405600D00077A045C0";
    attribute INIT_0D of inst : label is "72A04700D00076004780730051C0770051C072004780D00076A0470073405120";
    attribute INIT_0E of inst : label is "D00074405600722052C07770508073204680D000754047E07290525077405120";
    attribute INIT_0F of inst : label is "47E070F05360776054F073E04500D00070205600719053207780544073A045C0";
    attribute INIT_10 of inst : label is "537076C0562072005040D00071C047A0704053807720559072005420D0007100";
    attribute INIT_11 of inst : label is "570073804200D000730046A0752053407650569073E04140D000728047207480";
    attribute INIT_12 of inst : label is "4320D00073E045407650529075205740730042A0D0007380460075C0530075C0";
    attribute INIT_13 of inst : label is "72005020772051907040578071C043A0D0007200544076C05220748057707280";
    attribute INIT_14 of inst : label is "778050407190572070205200D00073E04100776050F070F05760710043E0D000";
    attribute INIT_15 of inst : label is "72905650754043E0D0007320428077705480722056C074405200D00073A041C0";
    attribute INIT_16 of inst : label is "3180E8DE06005460C84E02004060E8D5F80EC845F809D00072A0430077405520";
    attribute INIT_17 of inst : label is "06C046C0C86902C032C0E8F007404640C86003403240E8E707C04580C85703C0";
    attribute INIT_18 of inst : label is "C88400604200E90B058047C0C87B018033C0E90206404740C87202403340E8F9";
    attribute INIT_19 of inst : label is "C89F058033C0E92600605600C89604604200E91DFE08C88DF908E91404605600";
    attribute INIT_1A of inst : label is "3240E94102C046C0C8B106C032C0E93802404740C8A806403340E92F018047C0";
    attribute INIT_1B of inst : label is "02005460C8CC06004060E95303C04580C8C307C03180E94A03404640C8BA0740";
    attribute INIT_1C of inst : label is "F871F901C9D702003480F871FD70F87502003180C9D70000700001A0A080E95C";
    attribute INIT_1D of inst : label is "3E281200D000F578F577F177F178F173F573D000030034C0F770F87570001300";
    attribute INIT_1E of inst : label is "630003805480FD090700558007005180F9090380508005805600B4AB957F6954";
    attribute INIT_1F of inst : label is "45C006D055D00730513001E04240037050D005505620F20BF60B04C0670004C0";
    attribute INIT_20 of inst : label is "4260035051300510564002C04260034045C004786710050862E8038054200240";
    attribute INIT_21 of inst : label is "42800340456004286718055062D003905030026045A006B05610074050E001A0";
    attribute INIT_22 of inst : label is "62A803805080028045400670565007505090014042800340518004E0566002A0";
    attribute INIT_23 of inst : label is "569007505040010042A0031051D004A05670024042C003804500002867180598";
    attribute INIT_24 of inst : label is "02E0522004605680F30A038044A00070671005D06278036050E002A045000630";
    attribute INIT_25 of inst : label is "03A0444000C06700061062480350513002C044C005F056C00760542000C042C0";
    attribute INIT_26 of inst : label is "0330519002C044A005A056E007505470008042C002A052600420568001A04320";
    attribute INIT_27 of inst : label is "074054C0004042C0026052A0002056800160436003A04000011066E806506210";
    attribute INIT_28 of inst : label is "006056800120436003804060015866C8068061D8031051D002C0444005605710";
    attribute INIT_29 of inst : label is "019866A806A8619802E0522002C040000510573007305510000042C0022052E0";
    attribute INIT_2A of inst : label is "73805480FD797700558077005180F979738050800580560000C04380038040C0";
    attribute INIT_2B of inst : label is "FB70D000F602F872F906FE70F672F272FA70D0000220708074C0670074C06300";
    attribute INIT_2C of inst : label is "FB70EB58FF06F872FB70EB0AF077F575F570F571F003F077F575F570F571F073";
    attribute INIT_2D of inst : label is "FB70D000F803F700F077F705F872FB70F806F872EB0AF076F676F670F672F072";
    attribute INIT_2E of inst : label is "FF70F006F872FB06F872EB71F300F872F700FB70EB09F670F072F606F670F872";
    attribute INIT_2F of inst : label is "FB70EB58FF70FB00D000F003F773F777F003FB70EB36F072F672F200D000F802";
    attribute INIT_30 of inst : label is "F876F770F872FB70D000F803F876FF70F872FB70EB36FF72FB70EB71F272F672";
    attribute INIT_31 of inst : label is "EB59F773F001F876F770F872FB70EB59F672F202F076F676FE70F872FB70EADC";
    attribute INIT_32 of inst : label is "F872F370F876F370F872D000F072F670F076F670F072F601FE70F906FA73F200";
    attribute INIT_33 of inst : label is "F272FF70FB00EB37FB71FF71FB00D000FF01FB70F872FF70FB00EAEDFB00EB37";
    attribute INIT_34 of inst : label is "FF76F872FB00D000FE02F676F802F276FA70F002EB72FF72F806FB72EB36F672";
    attribute INIT_35 of inst : label is "F300F876FF70F872FB00D000F002F872F770F876F770F872FB00EAEFFB01EB58";
    attribute INIT_36 of inst : label is "FB00D000FF03FB70F876F770F872F300EB71F300F872F770FB00D000F702F872";
    attribute INIT_37 of inst : label is "CB53CB51CB06CB0AEB70F370F876F300F802EB5CFB70CB77D000F002FF70F872";
    attribute INIT_38 of inst : label is "CAEBCAE6CADFCAD8CAD6CACFCACBCABFCAB7CB77CB75CB6FCB68CB2BCB63CB5B";
    attribute INIT_39 of inst : label is "CB46CB42CB3DCB39CB33CB31CB2BCB19CB11CB0CCB06CB03CAFFCAFCCAF6CAF2";
    attribute INIT_3A of inst : label is "72FF92FF700096FF77FF9000700092FF73FF9000000070000000A080CB74CB4D";
    attribute INIT_3B of inst : label is "76FF96FF0000700003FFA37F72FF96FF720081FE7600920077FE87FE72008600";
    attribute INIT_3C of inst : label is "F900F0DB0000700001F4A1FC76FF92FF7600860073FE87FE72009200760081FE";
    attribute INIT_3D of inst : label is "F900F05BF900F06FF900F07BF900F08FF900F09BF900F0AFF900F0BBF900F0CF";
    attribute INIT_3E of inst : label is "CAD6CB0ACAF6CB03CAB7CABF00007000115EA0E4D000F02FF900F03BF900F04F";
    attribute INIT_3F of inst : label is "EADFCB03CAEBCB2BCAB7CB19CAD6EBEF00007000119AA0C0EB19CB06CB19CB19";
  begin
  inst : RAMB16_S9
      --pragma translate_off
      generic map (
        INITP_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
        INITP_07 => x"0000000000000000000000000000000000000000000000000000000000000000",

        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 0),
        DOP  => open,
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "00000000",
        DIP  => "0",
        EN   => '1',
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
